entity renormalizer_tb is
end renormalizer_tb;

architecture behave of renormalizer_tb is
begin
end behave;
