entity renormalizer is
end renormalizer;

architecture behave of renormalizer is 
begin
end behave;